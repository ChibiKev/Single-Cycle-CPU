library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_Control_vlg_vec_tst is
end Chen_Kevin_Control_vlg_vec_tst;
