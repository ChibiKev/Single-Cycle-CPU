Library ieee;
use ieee.std_logic_1164.all;

entity Chen_Kevin_Bitwise_NOT is
port(
			Chen_Kevin_a: in std_logic_vector(31 downto 0);
			Chen_Kevin_result: out std_logic_vector(31 downto 0)
			);
end Chen_Kevin_Bitwise_NOT;

architecture arch of Chen_Kevin_Bitwise_NOT is

begin
			Chen_Kevin_result <= NOT Chen_Kevin_a;
end arch;