library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_Single_Cycle_CPU_Board is
    port(
        Chen_Kevin_Segment_A0: out    vl_logic;
        Chen_Kevin_Clock: in     vl_logic;
        Chen_Keivn_Reset: in     vl_logic;
        Chen_Kevin_Segment_B0: out    vl_logic;
        Chen_Kevin_Segment_C0: out    vl_logic;
        Chen_Kevin_Segment_D0: out    vl_logic;
        Chen_Kevin_Segment_E0: out    vl_logic;
        Chen_Kevin_Segment_F0: out    vl_logic;
        Chen_Kevin_Segment_G0: out    vl_logic;
        Chen_Kevin_Segment_A1: out    vl_logic;
        Chen_Kevin_Segment_B1: out    vl_logic;
        Chen_Kevin_Segment_C1: out    vl_logic;
        Chen_Kevin_Segment_D1: out    vl_logic;
        Chen_Kevin_Segment_E1: out    vl_logic;
        Chen_Kevin_Segment_F1: out    vl_logic;
        Chen_Kevin_Segment_G1: out    vl_logic;
        Chen_Kevin_Segment_A2: out    vl_logic;
        Chen_Kevin_Segment_B2: out    vl_logic;
        Chen_Kevin_Segment_C2: out    vl_logic;
        Chen_Kevin_Segment_D2: out    vl_logic;
        Chen_Kevin_Segment_E2: out    vl_logic;
        Chen_Kevin_Segment_F2: out    vl_logic;
        Chen_Kevin_Segment_G2: out    vl_logic;
        Chen_Kevin_Segment_A3: out    vl_logic;
        Chen_Kevin_Segment_B3: out    vl_logic;
        Chen_Kevin_Segment_C3: out    vl_logic;
        Chen_Kevin_Segment_D3: out    vl_logic;
        Chen_Kevin_Segment_E3: out    vl_logic;
        Chen_Kevin_Segment_F3: out    vl_logic;
        Chen_Kevin_Segment_G3: out    vl_logic;
        Chen_Kevin_Segment_A4: out    vl_logic;
        Chen_Kevin_Segment_B4: out    vl_logic;
        Chen_Kevin_Segment_C4: out    vl_logic;
        Chen_Kevin_Segment_D4: out    vl_logic;
        Chen_Kevin_Segment_E4: out    vl_logic;
        Chen_Kevin_Segment_F4: out    vl_logic;
        Chen_Kevin_Segment_G4: out    vl_logic;
        Chen_Kevin_Segment_A5: out    vl_logic;
        Chen_Kevin_Segment_B5: out    vl_logic;
        Chen_Kevin_Segment_C5: out    vl_logic;
        Chen_Kevin_Segment_D5: out    vl_logic;
        Chen_Kevin_Segment_E5: out    vl_logic;
        Chen_Kevin_Segment_F5: out    vl_logic;
        Chen_Kevin_Segment_G5: out    vl_logic;
        Chen_Kevin_Segment_A6: out    vl_logic;
        Chen_Kevin_Segment_B6: out    vl_logic;
        Chen_Kevin_Segment_C6: out    vl_logic;
        Chen_Kevin_Segment_D6: out    vl_logic;
        Chen_Kevin_Segment_E6: out    vl_logic;
        Chen_Kevin_Segment_F6: out    vl_logic;
        Chen_Kevin_Segment_G6: out    vl_logic;
        Chen_Kevin_Segment_A7: out    vl_logic;
        Chen_Kevin_Segment_B7: out    vl_logic;
        Chen_Kevin_Segment_C7: out    vl_logic;
        Chen_Kevin_Segment_D7: out    vl_logic;
        Chen_Kevin_Segment_E7: out    vl_logic;
        Chen_Kevin_Segment_F7: out    vl_logic;
        Chen_Kevin_Segment_G7: out    vl_logic;
        Chen_Kevin_Op   : out    vl_logic_vector(3 downto 0)
    );
end Chen_Kevin_Single_Cycle_CPU_Board;
