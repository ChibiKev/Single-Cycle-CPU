library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_Add_By_Four_vlg_sample_tst is
    port(
        Chen_Kevin_a    : in     vl_logic_vector(31 downto 0);
        sampler_tx      : out    vl_logic
    );
end Chen_Kevin_Add_By_Four_vlg_sample_tst;
