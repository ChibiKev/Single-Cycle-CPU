library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_Single_Cycle_CPU_Board_vlg_check_tst is
    port(
        Chen_Kevin_Op   : in     vl_logic_vector(3 downto 0);
        Chen_Kevin_Segment_A0: in     vl_logic;
        Chen_Kevin_Segment_A1: in     vl_logic;
        Chen_Kevin_Segment_A2: in     vl_logic;
        Chen_Kevin_Segment_A3: in     vl_logic;
        Chen_Kevin_Segment_A4: in     vl_logic;
        Chen_Kevin_Segment_A5: in     vl_logic;
        Chen_Kevin_Segment_A6: in     vl_logic;
        Chen_Kevin_Segment_A7: in     vl_logic;
        Chen_Kevin_Segment_B0: in     vl_logic;
        Chen_Kevin_Segment_B1: in     vl_logic;
        Chen_Kevin_Segment_B2: in     vl_logic;
        Chen_Kevin_Segment_B3: in     vl_logic;
        Chen_Kevin_Segment_B4: in     vl_logic;
        Chen_Kevin_Segment_B5: in     vl_logic;
        Chen_Kevin_Segment_B6: in     vl_logic;
        Chen_Kevin_Segment_B7: in     vl_logic;
        Chen_Kevin_Segment_C0: in     vl_logic;
        Chen_Kevin_Segment_C1: in     vl_logic;
        Chen_Kevin_Segment_C2: in     vl_logic;
        Chen_Kevin_Segment_C3: in     vl_logic;
        Chen_Kevin_Segment_C4: in     vl_logic;
        Chen_Kevin_Segment_C5: in     vl_logic;
        Chen_Kevin_Segment_C6: in     vl_logic;
        Chen_Kevin_Segment_C7: in     vl_logic;
        Chen_Kevin_Segment_D0: in     vl_logic;
        Chen_Kevin_Segment_D1: in     vl_logic;
        Chen_Kevin_Segment_D2: in     vl_logic;
        Chen_Kevin_Segment_D3: in     vl_logic;
        Chen_Kevin_Segment_D4: in     vl_logic;
        Chen_Kevin_Segment_D5: in     vl_logic;
        Chen_Kevin_Segment_D6: in     vl_logic;
        Chen_Kevin_Segment_D7: in     vl_logic;
        Chen_Kevin_Segment_E0: in     vl_logic;
        Chen_Kevin_Segment_E1: in     vl_logic;
        Chen_Kevin_Segment_E2: in     vl_logic;
        Chen_Kevin_Segment_E3: in     vl_logic;
        Chen_Kevin_Segment_E4: in     vl_logic;
        Chen_Kevin_Segment_E5: in     vl_logic;
        Chen_Kevin_Segment_E6: in     vl_logic;
        Chen_Kevin_Segment_E7: in     vl_logic;
        Chen_Kevin_Segment_F0: in     vl_logic;
        Chen_Kevin_Segment_F1: in     vl_logic;
        Chen_Kevin_Segment_F2: in     vl_logic;
        Chen_Kevin_Segment_F3: in     vl_logic;
        Chen_Kevin_Segment_F4: in     vl_logic;
        Chen_Kevin_Segment_F5: in     vl_logic;
        Chen_Kevin_Segment_F6: in     vl_logic;
        Chen_Kevin_Segment_F7: in     vl_logic;
        Chen_Kevin_Segment_G0: in     vl_logic;
        Chen_Kevin_Segment_G1: in     vl_logic;
        Chen_Kevin_Segment_G2: in     vl_logic;
        Chen_Kevin_Segment_G3: in     vl_logic;
        Chen_Kevin_Segment_G4: in     vl_logic;
        Chen_Kevin_Segment_G5: in     vl_logic;
        Chen_Kevin_Segment_G6: in     vl_logic;
        Chen_Kevin_Segment_G7: in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Chen_Kevin_Single_Cycle_CPU_Board_vlg_check_tst;
