library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;  

entity Chen_Kevin_Instruction is
port (
 Chen_Kevin_Read_Address: in std_logic_vector(31 downto 0);
 Chen_Kevin_Instruction: out  std_logic_vector(31 downto 0)
);
end Chen_Kevin_Instruction;

architecture arch of Chen_Kevin_Instruction is
signal Chen_Kevin_ROM_Address: std_logic_vector(4 downto 0);
 type Chen_Kevin_ROM_Type is array (0 to 31 ) of std_logic_vector(31 downto 0);
 constant Chen_Kevin_ROM_Data: Chen_Kevin_ROM_Type:=(
   "10101101000100000000000000000000",
	--101011 sw | 01000 register 8, $t0 | 10000 register 16, $s0. $t0 = $s0
   "00000001000100010100000000000010", 
	--000000 R-Type | 01000 $t0 | 10001 $s1 | 01000 $t0 | 00000 | 000010 add. $t0 += $s1
   "00000001000100010100000000000010", 
	--000000 R-Type | 01000 $t0 | 10001 $s1 | 01000 $t0 | 00000 | 000010 add. $t0 += $s1
   "00000001000100010100000000000010", 
	--000000 R-Type | 01000 $t0 | 10001 $s1 | 01000 $t0 | 00000 | 000010 add. $t0 += $s1
   "00000001000100100100000000000011", 
	--000000 R-Type | 01000 $t0 | 10010 $s2 | 01000 $t0 | 00000 | 000011 sub. $t0 -= $s2
   "00000000000000000000000000000000", 
   "00000000000000000000000000000000", 
   "00000000000000000000000000000000", 
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000"
  );
begin

 Chen_Kevin_ROM_Address <= Chen_Kevin_Read_Address(5 downto 1);
  Chen_Kevin_Instruction <= Chen_Kevin_ROM_Data((to_integer(unsigned(Chen_Kevin_ROM_Address)))/2) when Chen_Kevin_Read_Address < x"00000020" else x"00000000";

end arch;